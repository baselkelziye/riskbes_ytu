module partial_product (
 input  [31:0] muler_i, mulcand_i,
 output [31:0] pp0_o,  pp1_o,  pp2_o,  pp3_o,  pp4_o,  pp5_o,  pp6_o,  pp7_o, 
               pp8_o,  pp9_o,  pp10_o, pp11_o, pp12_o, pp13_o, pp14_o, pp15_o,
               pp16_o, pp17_o, pp18_o, pp19_o, pp20_o, pp21_o, pp22_o, pp23_o,
               pp24_o, pp25_o, pp26_o, pp27_o, pp28_o, pp29_o, pp30_o, pp31_o
);
   assign pp0_o[0]   = muler_i[0]  & mulcand_i[0];
   assign pp1_o[0]   = muler_i[0]  & mulcand_i[1];
   assign pp2_o[0]   = muler_i[0]  & mulcand_i[2];
   assign pp3_o[0]   = muler_i[0]  & mulcand_i[3];
   assign pp4_o[0]   = muler_i[0]  & mulcand_i[4];
   assign pp5_o[0]   = muler_i[0]  & mulcand_i[5];
   assign pp6_o[0]   = muler_i[0]  & mulcand_i[6];
   assign pp7_o[0]   = muler_i[0]  & mulcand_i[7];
   assign pp8_o[0]   = muler_i[0]  & mulcand_i[8];
   assign pp9_o[0]   = muler_i[0]  & mulcand_i[9];
   assign pp10_o[0]  = muler_i[0]  & mulcand_i[10];
   assign pp11_o[0]  = muler_i[0]  & mulcand_i[11];
   assign pp12_o[0]  = muler_i[0]  & mulcand_i[12];
   assign pp13_o[0]  = muler_i[0]  & mulcand_i[13];
   assign pp14_o[0]  = muler_i[0]  & mulcand_i[14];
   assign pp15_o[0]  = muler_i[0]  & mulcand_i[15];
   assign pp16_o[0]  = muler_i[0]  & mulcand_i[16];
   assign pp17_o[0]  = muler_i[0]  & mulcand_i[17];
   assign pp18_o[0]  = muler_i[0]  & mulcand_i[18];
   assign pp19_o[0]  = muler_i[0]  & mulcand_i[19];
   assign pp20_o[0]  = muler_i[0]  & mulcand_i[20];
   assign pp21_o[0]  = muler_i[0]  & mulcand_i[21];
   assign pp22_o[0]  = muler_i[0]  & mulcand_i[22];
   assign pp23_o[0]  = muler_i[0]  & mulcand_i[23];
   assign pp24_o[0]  = muler_i[0]  & mulcand_i[24];
   assign pp25_o[0]  = muler_i[0]  & mulcand_i[25];
   assign pp26_o[0]  = muler_i[0]  & mulcand_i[26];
   assign pp27_o[0]  = muler_i[0]  & mulcand_i[27];
   assign pp28_o[0]  = muler_i[0]  & mulcand_i[28];
   assign pp29_o[0]  = muler_i[0]  & mulcand_i[29];
   assign pp30_o[0]  = muler_i[0]  & mulcand_i[30];
   assign pp31_o[0]  = muler_i[0]  & mulcand_i[31];

   assign pp0_o[1]   = muler_i[1]  & mulcand_i[0];
   assign pp1_o[1]   = muler_i[1]  & mulcand_i[1];
   assign pp2_o[1]   = muler_i[1]  & mulcand_i[2];
   assign pp3_o[1]   = muler_i[1]  & mulcand_i[3];
   assign pp4_o[1]   = muler_i[1]  & mulcand_i[4];
   assign pp5_o[1]   = muler_i[1]  & mulcand_i[5];
   assign pp6_o[1]   = muler_i[1]  & mulcand_i[6];
   assign pp7_o[1]   = muler_i[1]  & mulcand_i[7];
   assign pp8_o[1]   = muler_i[1]  & mulcand_i[8];
   assign pp9_o[1]   = muler_i[1]  & mulcand_i[9];
   assign pp10_o[1]  = muler_i[1]  & mulcand_i[10];
   assign pp11_o[1]  = muler_i[1]  & mulcand_i[11];
   assign pp12_o[1]  = muler_i[1]  & mulcand_i[12];
   assign pp13_o[1]  = muler_i[1]  & mulcand_i[13];
   assign pp14_o[1]  = muler_i[1]  & mulcand_i[14];
   assign pp15_o[1]  = muler_i[1]  & mulcand_i[15];
   assign pp16_o[1]  = muler_i[1]  & mulcand_i[16];
   assign pp17_o[1]  = muler_i[1]  & mulcand_i[17];
   assign pp18_o[1]  = muler_i[1]  & mulcand_i[18];
   assign pp19_o[1]  = muler_i[1]  & mulcand_i[19];
   assign pp20_o[1]  = muler_i[1]  & mulcand_i[20];
   assign pp21_o[1]  = muler_i[1]  & mulcand_i[21];
   assign pp22_o[1]  = muler_i[1]  & mulcand_i[22];
   assign pp23_o[1]  = muler_i[1]  & mulcand_i[23];
   assign pp24_o[1]  = muler_i[1]  & mulcand_i[24];
   assign pp25_o[1]  = muler_i[1]  & mulcand_i[25];
   assign pp26_o[1]  = muler_i[1]  & mulcand_i[26];
   assign pp27_o[1]  = muler_i[1]  & mulcand_i[27];
   assign pp28_o[1]  = muler_i[1]  & mulcand_i[28];
   assign pp29_o[1]  = muler_i[1]  & mulcand_i[29];
   assign pp30_o[1]  = muler_i[1]  & mulcand_i[30];
   assign pp31_o[1]  = muler_i[1]  & mulcand_i[31];

   assign pp0_o[2]   = muler_i[2]  & mulcand_i[0];
   assign pp1_o[2]   = muler_i[2]  & mulcand_i[1];
   assign pp2_o[2]   = muler_i[2]  & mulcand_i[2];
   assign pp3_o[2]   = muler_i[2]  & mulcand_i[3];
   assign pp4_o[2]   = muler_i[2]  & mulcand_i[4];
   assign pp5_o[2]   = muler_i[2]  & mulcand_i[5];
   assign pp6_o[2]   = muler_i[2]  & mulcand_i[6];
   assign pp7_o[2]   = muler_i[2]  & mulcand_i[7];
   assign pp8_o[2]   = muler_i[2]  & mulcand_i[8];
   assign pp9_o[2]   = muler_i[2]  & mulcand_i[9];
   assign pp10_o[2]  = muler_i[2]  & mulcand_i[10];
   assign pp11_o[2]  = muler_i[2]  & mulcand_i[11];
   assign pp12_o[2]  = muler_i[2]  & mulcand_i[12];
   assign pp13_o[2]  = muler_i[2]  & mulcand_i[13];
   assign pp14_o[2]  = muler_i[2]  & mulcand_i[14];
   assign pp15_o[2]  = muler_i[2]  & mulcand_i[15];
   assign pp16_o[2]  = muler_i[2]  & mulcand_i[16];
   assign pp17_o[2]  = muler_i[2]  & mulcand_i[17];
   assign pp18_o[2]  = muler_i[2]  & mulcand_i[18];
   assign pp19_o[2]  = muler_i[2]  & mulcand_i[19];
   assign pp20_o[2]  = muler_i[2]  & mulcand_i[20];
   assign pp21_o[2]  = muler_i[2]  & mulcand_i[21];
   assign pp22_o[2]  = muler_i[2]  & mulcand_i[22];
   assign pp23_o[2]  = muler_i[2]  & mulcand_i[23];
   assign pp24_o[2]  = muler_i[2]  & mulcand_i[24];
   assign pp25_o[2]  = muler_i[2]  & mulcand_i[25];
   assign pp26_o[2]  = muler_i[2]  & mulcand_i[26];
   assign pp27_o[2]  = muler_i[2]  & mulcand_i[27];
   assign pp28_o[2]  = muler_i[2]  & mulcand_i[28];
   assign pp29_o[2]  = muler_i[2]  & mulcand_i[29];
   assign pp30_o[2]  = muler_i[2]  & mulcand_i[30];
   assign pp31_o[2]  = muler_i[2]  & mulcand_i[31];

   assign pp0_o[3]   = muler_i[3]  & mulcand_i[0];
   assign pp1_o[3]   = muler_i[3]  & mulcand_i[1];
   assign pp2_o[3]   = muler_i[3]  & mulcand_i[2];
   assign pp3_o[3]   = muler_i[3]  & mulcand_i[3];
   assign pp4_o[3]   = muler_i[3]  & mulcand_i[4];
   assign pp5_o[3]   = muler_i[3]  & mulcand_i[5];
   assign pp6_o[3]   = muler_i[3]  & mulcand_i[6];
   assign pp7_o[3]   = muler_i[3]  & mulcand_i[7];
   assign pp8_o[3]   = muler_i[3]  & mulcand_i[8];
   assign pp9_o[3]   = muler_i[3]  & mulcand_i[9];
   assign pp10_o[3]  = muler_i[3]  & mulcand_i[10];
   assign pp11_o[3]  = muler_i[3]  & mulcand_i[11];
   assign pp12_o[3]  = muler_i[3]  & mulcand_i[12];
   assign pp13_o[3]  = muler_i[3]  & mulcand_i[13];
   assign pp14_o[3]  = muler_i[3]  & mulcand_i[14];
   assign pp15_o[3]  = muler_i[3]  & mulcand_i[15];
   assign pp16_o[3]  = muler_i[3]  & mulcand_i[16];
   assign pp17_o[3]  = muler_i[3]  & mulcand_i[17];
   assign pp18_o[3]  = muler_i[3]  & mulcand_i[18];
   assign pp19_o[3]  = muler_i[3]  & mulcand_i[19];
   assign pp20_o[3]  = muler_i[3]  & mulcand_i[20];
   assign pp21_o[3]  = muler_i[3]  & mulcand_i[21];
   assign pp22_o[3]  = muler_i[3]  & mulcand_i[22];
   assign pp23_o[3]  = muler_i[3]  & mulcand_i[23];
   assign pp24_o[3]  = muler_i[3]  & mulcand_i[24];
   assign pp25_o[3]  = muler_i[3]  & mulcand_i[25];
   assign pp26_o[3]  = muler_i[3]  & mulcand_i[26];
   assign pp27_o[3]  = muler_i[3]  & mulcand_i[27];
   assign pp28_o[3]  = muler_i[3]  & mulcand_i[28];
   assign pp29_o[3]  = muler_i[3]  & mulcand_i[29];
   assign pp30_o[3]  = muler_i[3]  & mulcand_i[30];
   assign pp31_o[3]  = muler_i[3]  & mulcand_i[31];

   assign pp0_o[4]   = muler_i[4]  & mulcand_i[0];
   assign pp1_o[4]   = muler_i[4]  & mulcand_i[1];
   assign pp2_o[4]   = muler_i[4]  & mulcand_i[2];
   assign pp3_o[4]   = muler_i[4]  & mulcand_i[3];
   assign pp4_o[4]   = muler_i[4]  & mulcand_i[4];
   assign pp5_o[4]   = muler_i[4]  & mulcand_i[5];
   assign pp6_o[4]   = muler_i[4]  & mulcand_i[6];
   assign pp7_o[4]   = muler_i[4]  & mulcand_i[7];
   assign pp8_o[4]   = muler_i[4]  & mulcand_i[8];
   assign pp9_o[4]   = muler_i[4]  & mulcand_i[9];
   assign pp10_o[4]  = muler_i[4]  & mulcand_i[10];
   assign pp11_o[4]  = muler_i[4]  & mulcand_i[11];
   assign pp12_o[4]  = muler_i[4]  & mulcand_i[12];
   assign pp13_o[4]  = muler_i[4]  & mulcand_i[13];
   assign pp14_o[4]  = muler_i[4]  & mulcand_i[14];
   assign pp15_o[4]  = muler_i[4]  & mulcand_i[15];
   assign pp16_o[4]  = muler_i[4]  & mulcand_i[16];
   assign pp17_o[4]  = muler_i[4]  & mulcand_i[17];
   assign pp18_o[4]  = muler_i[4]  & mulcand_i[18];
   assign pp19_o[4]  = muler_i[4]  & mulcand_i[19];
   assign pp20_o[4]  = muler_i[4]  & mulcand_i[20];
   assign pp21_o[4]  = muler_i[4]  & mulcand_i[21];
   assign pp22_o[4]  = muler_i[4]  & mulcand_i[22];
   assign pp23_o[4]  = muler_i[4]  & mulcand_i[23];
   assign pp24_o[4]  = muler_i[4]  & mulcand_i[24];
   assign pp25_o[4]  = muler_i[4]  & mulcand_i[25];
   assign pp26_o[4]  = muler_i[4]  & mulcand_i[26];
   assign pp27_o[4]  = muler_i[4]  & mulcand_i[27];
   assign pp28_o[4]  = muler_i[4]  & mulcand_i[28];
   assign pp29_o[4]  = muler_i[4]  & mulcand_i[29];
   assign pp30_o[4]  = muler_i[4]  & mulcand_i[30];
   assign pp31_o[4]  = muler_i[4]  & mulcand_i[31];

   assign pp0_o[5]   = muler_i[5]  & mulcand_i[0];
   assign pp1_o[5]   = muler_i[5]  & mulcand_i[1];
   assign pp2_o[5]   = muler_i[5]  & mulcand_i[2];
   assign pp3_o[5]   = muler_i[5]  & mulcand_i[3];
   assign pp4_o[5]   = muler_i[5]  & mulcand_i[4];
   assign pp5_o[5]   = muler_i[5]  & mulcand_i[5];
   assign pp6_o[5]   = muler_i[5]  & mulcand_i[6];
   assign pp7_o[5]   = muler_i[5]  & mulcand_i[7];
   assign pp8_o[5]   = muler_i[5]  & mulcand_i[8];
   assign pp9_o[5]   = muler_i[5]  & mulcand_i[9];
   assign pp10_o[5]  = muler_i[5]  & mulcand_i[10];
   assign pp11_o[5]  = muler_i[5]  & mulcand_i[11];
   assign pp12_o[5]  = muler_i[5]  & mulcand_i[12];
   assign pp13_o[5]  = muler_i[5]  & mulcand_i[13];
   assign pp14_o[5]  = muler_i[5]  & mulcand_i[14];
   assign pp15_o[5]  = muler_i[5]  & mulcand_i[15];
   assign pp16_o[5]  = muler_i[5]  & mulcand_i[16];
   assign pp17_o[5]  = muler_i[5]  & mulcand_i[17];
   assign pp18_o[5]  = muler_i[5]  & mulcand_i[18];
   assign pp19_o[5]  = muler_i[5]  & mulcand_i[19];
   assign pp20_o[5]  = muler_i[5]  & mulcand_i[20];
   assign pp21_o[5]  = muler_i[5]  & mulcand_i[21];
   assign pp22_o[5]  = muler_i[5]  & mulcand_i[22];
   assign pp23_o[5]  = muler_i[5]  & mulcand_i[23];
   assign pp24_o[5]  = muler_i[5]  & mulcand_i[24];
   assign pp25_o[5]  = muler_i[5]  & mulcand_i[25];
   assign pp26_o[5]  = muler_i[5]  & mulcand_i[26];
   assign pp27_o[5]  = muler_i[5]  & mulcand_i[27];
   assign pp28_o[5]  = muler_i[5]  & mulcand_i[28];
   assign pp29_o[5]  = muler_i[5]  & mulcand_i[29];
   assign pp30_o[5]  = muler_i[5]  & mulcand_i[30];
   assign pp31_o[5]  = muler_i[5]  & mulcand_i[31];

   assign pp0_o[6]   = muler_i[6]  & mulcand_i[0];
   assign pp1_o[6]   = muler_i[6]  & mulcand_i[1];
   assign pp2_o[6]   = muler_i[6]  & mulcand_i[2];
   assign pp3_o[6]   = muler_i[6]  & mulcand_i[3];
   assign pp4_o[6]   = muler_i[6]  & mulcand_i[4];
   assign pp5_o[6]   = muler_i[6]  & mulcand_i[5];
   assign pp6_o[6]   = muler_i[6]  & mulcand_i[6];
   assign pp7_o[6]   = muler_i[6]  & mulcand_i[7];
   assign pp8_o[6]   = muler_i[6]  & mulcand_i[8];
   assign pp9_o[6]   = muler_i[6]  & mulcand_i[9];
   assign pp10_o[6]  = muler_i[6]  & mulcand_i[10];
   assign pp11_o[6]  = muler_i[6]  & mulcand_i[11];
   assign pp12_o[6]  = muler_i[6]  & mulcand_i[12];
   assign pp13_o[6]  = muler_i[6]  & mulcand_i[13];
   assign pp14_o[6]  = muler_i[6]  & mulcand_i[14];
   assign pp15_o[6]  = muler_i[6]  & mulcand_i[15];
   assign pp16_o[6]  = muler_i[6]  & mulcand_i[16];
   assign pp17_o[6]  = muler_i[6]  & mulcand_i[17];
   assign pp18_o[6]  = muler_i[6]  & mulcand_i[18];
   assign pp19_o[6]  = muler_i[6]  & mulcand_i[19];
   assign pp20_o[6]  = muler_i[6]  & mulcand_i[20];
   assign pp21_o[6]  = muler_i[6]  & mulcand_i[21];
   assign pp22_o[6]  = muler_i[6]  & mulcand_i[22];
   assign pp23_o[6]  = muler_i[6]  & mulcand_i[23];
   assign pp24_o[6]  = muler_i[6]  & mulcand_i[24];
   assign pp25_o[6]  = muler_i[6]  & mulcand_i[25];
   assign pp26_o[6]  = muler_i[6]  & mulcand_i[26];
   assign pp27_o[6]  = muler_i[6]  & mulcand_i[27];
   assign pp28_o[6]  = muler_i[6]  & mulcand_i[28];
   assign pp29_o[6]  = muler_i[6]  & mulcand_i[29];
   assign pp30_o[6]  = muler_i[6]  & mulcand_i[30];
   assign pp31_o[6]  = muler_i[6]  & mulcand_i[31];

   assign pp0_o[7]   = muler_i[7]  & mulcand_i[0];
   assign pp1_o[7]   = muler_i[7]  & mulcand_i[1];
   assign pp2_o[7]   = muler_i[7]  & mulcand_i[2];
   assign pp3_o[7]   = muler_i[7]  & mulcand_i[3];
   assign pp4_o[7]   = muler_i[7]  & mulcand_i[4];
   assign pp5_o[7]   = muler_i[7]  & mulcand_i[5];
   assign pp6_o[7]   = muler_i[7]  & mulcand_i[6];
   assign pp7_o[7]   = muler_i[7]  & mulcand_i[7];
   assign pp8_o[7]   = muler_i[7]  & mulcand_i[8];
   assign pp9_o[7]   = muler_i[7]  & mulcand_i[9];
   assign pp10_o[7]  = muler_i[7]  & mulcand_i[10];
   assign pp11_o[7]  = muler_i[7]  & mulcand_i[11];
   assign pp12_o[7]  = muler_i[7]  & mulcand_i[12];
   assign pp13_o[7]  = muler_i[7]  & mulcand_i[13];
   assign pp14_o[7]  = muler_i[7]  & mulcand_i[14];
   assign pp15_o[7]  = muler_i[7]  & mulcand_i[15];
   assign pp16_o[7]  = muler_i[7]  & mulcand_i[16];
   assign pp17_o[7]  = muler_i[7]  & mulcand_i[17];
   assign pp18_o[7]  = muler_i[7]  & mulcand_i[18];
   assign pp19_o[7]  = muler_i[7]  & mulcand_i[19];
   assign pp20_o[7]  = muler_i[7]  & mulcand_i[20];
   assign pp21_o[7]  = muler_i[7]  & mulcand_i[21];
   assign pp22_o[7]  = muler_i[7]  & mulcand_i[22];
   assign pp23_o[7]  = muler_i[7]  & mulcand_i[23];
   assign pp24_o[7]  = muler_i[7]  & mulcand_i[24];
   assign pp25_o[7]  = muler_i[7]  & mulcand_i[25];
   assign pp26_o[7]  = muler_i[7]  & mulcand_i[26];
   assign pp27_o[7]  = muler_i[7]  & mulcand_i[27];
   assign pp28_o[7]  = muler_i[7]  & mulcand_i[28];
   assign pp29_o[7]  = muler_i[7]  & mulcand_i[29];
   assign pp30_o[7]  = muler_i[7]  & mulcand_i[30];
   assign pp31_o[7]  = muler_i[7]  & mulcand_i[31];

   assign pp0_o[8]   = muler_i[8]  & mulcand_i[0];
   assign pp1_o[8]   = muler_i[8]  & mulcand_i[1];
   assign pp2_o[8]   = muler_i[8]  & mulcand_i[2];
   assign pp3_o[8]   = muler_i[8]  & mulcand_i[3];
   assign pp4_o[8]   = muler_i[8]  & mulcand_i[4];
   assign pp5_o[8]   = muler_i[8]  & mulcand_i[5];
   assign pp6_o[8]   = muler_i[8]  & mulcand_i[6];
   assign pp7_o[8]   = muler_i[8]  & mulcand_i[7];
   assign pp8_o[8]   = muler_i[8]  & mulcand_i[8];
   assign pp9_o[8]   = muler_i[8]  & mulcand_i[9];
   assign pp10_o[8]  = muler_i[8]  & mulcand_i[10];
   assign pp11_o[8]  = muler_i[8]  & mulcand_i[11];
   assign pp12_o[8]  = muler_i[8]  & mulcand_i[12];
   assign pp13_o[8]  = muler_i[8]  & mulcand_i[13];
   assign pp14_o[8]  = muler_i[8]  & mulcand_i[14];
   assign pp15_o[8]  = muler_i[8]  & mulcand_i[15];
   assign pp16_o[8]  = muler_i[8]  & mulcand_i[16];
   assign pp17_o[8]  = muler_i[8]  & mulcand_i[17];
   assign pp18_o[8]  = muler_i[8]  & mulcand_i[18];
   assign pp19_o[8]  = muler_i[8]  & mulcand_i[19];
   assign pp20_o[8]  = muler_i[8]  & mulcand_i[20];
   assign pp21_o[8]  = muler_i[8]  & mulcand_i[21];
   assign pp22_o[8]  = muler_i[8]  & mulcand_i[22];
   assign pp23_o[8]  = muler_i[8]  & mulcand_i[23];
   assign pp24_o[8]  = muler_i[8]  & mulcand_i[24];
   assign pp25_o[8]  = muler_i[8]  & mulcand_i[25];
   assign pp26_o[8]  = muler_i[8]  & mulcand_i[26];
   assign pp27_o[8]  = muler_i[8]  & mulcand_i[27];
   assign pp28_o[8]  = muler_i[8]  & mulcand_i[28];
   assign pp29_o[8]  = muler_i[8]  & mulcand_i[29];
   assign pp30_o[8]  = muler_i[8]  & mulcand_i[30];
   assign pp31_o[8]  = muler_i[8]  & mulcand_i[31];

   assign pp0_o[9]   = muler_i[9]  & mulcand_i[0];
   assign pp1_o[9]   = muler_i[9]  & mulcand_i[1];
   assign pp2_o[9]   = muler_i[9]  & mulcand_i[2];
   assign pp3_o[9]   = muler_i[9]  & mulcand_i[3];
   assign pp4_o[9]   = muler_i[9]  & mulcand_i[4];
   assign pp5_o[9]   = muler_i[9]  & mulcand_i[5];
   assign pp6_o[9]   = muler_i[9]  & mulcand_i[6];
   assign pp7_o[9]   = muler_i[9]  & mulcand_i[7];
   assign pp8_o[9]   = muler_i[9]  & mulcand_i[8];
   assign pp9_o[9]   = muler_i[9]  & mulcand_i[9];
   assign pp10_o[9]  = muler_i[9]  & mulcand_i[10];
   assign pp11_o[9]  = muler_i[9]  & mulcand_i[11];
   assign pp12_o[9]  = muler_i[9]  & mulcand_i[12];
   assign pp13_o[9]  = muler_i[9]  & mulcand_i[13];
   assign pp14_o[9]  = muler_i[9]  & mulcand_i[14];
   assign pp15_o[9]  = muler_i[9]  & mulcand_i[15];
   assign pp16_o[9]  = muler_i[9]  & mulcand_i[16];
   assign pp17_o[9]  = muler_i[9]  & mulcand_i[17];
   assign pp18_o[9]  = muler_i[9]  & mulcand_i[18];
   assign pp19_o[9]  = muler_i[9]  & mulcand_i[19];
   assign pp20_o[9]  = muler_i[9]  & mulcand_i[20];
   assign pp21_o[9]  = muler_i[9]  & mulcand_i[21];
   assign pp22_o[9]  = muler_i[9]  & mulcand_i[22];
   assign pp23_o[9]  = muler_i[9]  & mulcand_i[23];
   assign pp24_o[9]  = muler_i[9]  & mulcand_i[24];
   assign pp25_o[9]  = muler_i[9]  & mulcand_i[25];
   assign pp26_o[9]  = muler_i[9]  & mulcand_i[26];
   assign pp27_o[9]  = muler_i[9]  & mulcand_i[27];
   assign pp28_o[9]  = muler_i[9]  & mulcand_i[28];
   assign pp29_o[9]  = muler_i[9]  & mulcand_i[29];
   assign pp30_o[9]  = muler_i[9]  & mulcand_i[30];
   assign pp31_o[9]  = muler_i[9]  & mulcand_i[31];

   assign pp0_o[10]  = muler_i[10] & mulcand_i[0];
   assign pp1_o[10]  = muler_i[10] & mulcand_i[1];
   assign pp2_o[10]  = muler_i[10] & mulcand_i[2];
   assign pp3_o[10]  = muler_i[10] & mulcand_i[3];
   assign pp4_o[10]  = muler_i[10] & mulcand_i[4];
   assign pp5_o[10]  = muler_i[10] & mulcand_i[5];
   assign pp6_o[10]  = muler_i[10] & mulcand_i[6];
   assign pp7_o[10]  = muler_i[10] & mulcand_i[7];
   assign pp8_o[10]  = muler_i[10] & mulcand_i[8];
   assign pp9_o[10]  = muler_i[10] & mulcand_i[9];
   assign pp10_o[10] = muler_i[10] & mulcand_i[10];
   assign pp11_o[10] = muler_i[10] & mulcand_i[11];
   assign pp12_o[10] = muler_i[10] & mulcand_i[12];
   assign pp13_o[10] = muler_i[10] & mulcand_i[13];
   assign pp14_o[10] = muler_i[10] & mulcand_i[14];
   assign pp15_o[10] = muler_i[10] & mulcand_i[15];
   assign pp16_o[10] = muler_i[10] & mulcand_i[16];
   assign pp17_o[10] = muler_i[10] & mulcand_i[17];
   assign pp18_o[10] = muler_i[10] & mulcand_i[18];
   assign pp19_o[10] = muler_i[10] & mulcand_i[19];
   assign pp20_o[10] = muler_i[10] & mulcand_i[20];
   assign pp21_o[10] = muler_i[10] & mulcand_i[21];
   assign pp22_o[10] = muler_i[10] & mulcand_i[22];
   assign pp23_o[10] = muler_i[10] & mulcand_i[23];
   assign pp24_o[10] = muler_i[10] & mulcand_i[24];
   assign pp25_o[10] = muler_i[10] & mulcand_i[25];
   assign pp26_o[10] = muler_i[10] & mulcand_i[26];
   assign pp27_o[10] = muler_i[10] & mulcand_i[27];
   assign pp28_o[10] = muler_i[10] & mulcand_i[28];
   assign pp29_o[10] = muler_i[10] & mulcand_i[29];
   assign pp30_o[10] = muler_i[10] & mulcand_i[30];
   assign pp31_o[10] = muler_i[10] & mulcand_i[31];

   assign pp0_o[11]  = muler_i[11] & mulcand_i[0];
   assign pp1_o[11]  = muler_i[11] & mulcand_i[1];
   assign pp2_o[11]  = muler_i[11] & mulcand_i[2];
   assign pp3_o[11]  = muler_i[11] & mulcand_i[3];
   assign pp4_o[11]  = muler_i[11] & mulcand_i[4];
   assign pp5_o[11]  = muler_i[11] & mulcand_i[5];
   assign pp6_o[11]  = muler_i[11] & mulcand_i[6];
   assign pp7_o[11]  = muler_i[11] & mulcand_i[7];
   assign pp8_o[11]  = muler_i[11] & mulcand_i[8];
   assign pp9_o[11]  = muler_i[11] & mulcand_i[9];
   assign pp10_o[11] = muler_i[11] & mulcand_i[10];
   assign pp11_o[11] = muler_i[11] & mulcand_i[11];
   assign pp12_o[11] = muler_i[11] & mulcand_i[12];
   assign pp13_o[11] = muler_i[11] & mulcand_i[13];
   assign pp14_o[11] = muler_i[11] & mulcand_i[14];
   assign pp15_o[11] = muler_i[11] & mulcand_i[15];
   assign pp16_o[11] = muler_i[11] & mulcand_i[16];
   assign pp17_o[11] = muler_i[11] & mulcand_i[17];
   assign pp18_o[11] = muler_i[11] & mulcand_i[18];
   assign pp19_o[11] = muler_i[11] & mulcand_i[19];
   assign pp20_o[11] = muler_i[11] & mulcand_i[20];
   assign pp21_o[11] = muler_i[11] & mulcand_i[21];
   assign pp22_o[11] = muler_i[11] & mulcand_i[22];
   assign pp23_o[11] = muler_i[11] & mulcand_i[23];
   assign pp24_o[11] = muler_i[11] & mulcand_i[24];
   assign pp25_o[11] = muler_i[11] & mulcand_i[25];
   assign pp26_o[11] = muler_i[11] & mulcand_i[26];
   assign pp27_o[11] = muler_i[11] & mulcand_i[27];
   assign pp28_o[11] = muler_i[11] & mulcand_i[28];
   assign pp29_o[11] = muler_i[11] & mulcand_i[29];
   assign pp30_o[11] = muler_i[11] & mulcand_i[30];
   assign pp31_o[11] = muler_i[11] & mulcand_i[31];

   assign pp0_o[12]  = muler_i[12] & mulcand_i[0];
   assign pp1_o[12]  = muler_i[12] & mulcand_i[1];
   assign pp2_o[12]  = muler_i[12] & mulcand_i[2];
   assign pp3_o[12]  = muler_i[12] & mulcand_i[3];
   assign pp4_o[12]  = muler_i[12] & mulcand_i[4];
   assign pp5_o[12]  = muler_i[12] & mulcand_i[5];
   assign pp6_o[12]  = muler_i[12] & mulcand_i[6];
   assign pp7_o[12]  = muler_i[12] & mulcand_i[7];
   assign pp8_o[12]  = muler_i[12] & mulcand_i[8];
   assign pp9_o[12]  = muler_i[12] & mulcand_i[9];
   assign pp10_o[12] = muler_i[12] & mulcand_i[10];
   assign pp11_o[12] = muler_i[12] & mulcand_i[11];
   assign pp12_o[12] = muler_i[12] & mulcand_i[12];
   assign pp13_o[12] = muler_i[12] & mulcand_i[13];
   assign pp14_o[12] = muler_i[12] & mulcand_i[14];
   assign pp15_o[12] = muler_i[12] & mulcand_i[15];
   assign pp16_o[12] = muler_i[12] & mulcand_i[16];
   assign pp17_o[12] = muler_i[12] & mulcand_i[17];
   assign pp18_o[12] = muler_i[12] & mulcand_i[18];
   assign pp19_o[12] = muler_i[12] & mulcand_i[19];
   assign pp20_o[12] = muler_i[12] & mulcand_i[20];
   assign pp21_o[12] = muler_i[12] & mulcand_i[21];
   assign pp22_o[12] = muler_i[12] & mulcand_i[22];
   assign pp23_o[12] = muler_i[12] & mulcand_i[23];
   assign pp24_o[12] = muler_i[12] & mulcand_i[24];
   assign pp25_o[12] = muler_i[12] & mulcand_i[25];
   assign pp26_o[12] = muler_i[12] & mulcand_i[26];
   assign pp27_o[12] = muler_i[12] & mulcand_i[27];
   assign pp28_o[12] = muler_i[12] & mulcand_i[28];
   assign pp29_o[12] = muler_i[12] & mulcand_i[29];
   assign pp30_o[12] = muler_i[12] & mulcand_i[30];
   assign pp31_o[12] = muler_i[12] & mulcand_i[31];

   assign pp0_o[13]  = muler_i[13] & mulcand_i[0];
   assign pp1_o[13]  = muler_i[13] & mulcand_i[1];
   assign pp2_o[13]  = muler_i[13] & mulcand_i[2];
   assign pp3_o[13]  = muler_i[13] & mulcand_i[3];
   assign pp4_o[13]  = muler_i[13] & mulcand_i[4];
   assign pp5_o[13]  = muler_i[13] & mulcand_i[5];
   assign pp6_o[13]  = muler_i[13] & mulcand_i[6];
   assign pp7_o[13]  = muler_i[13] & mulcand_i[7];
   assign pp8_o[13]  = muler_i[13] & mulcand_i[8];
   assign pp9_o[13]  = muler_i[13] & mulcand_i[9];
   assign pp10_o[13] = muler_i[13] & mulcand_i[10];
   assign pp11_o[13] = muler_i[13] & mulcand_i[11];
   assign pp12_o[13] = muler_i[13] & mulcand_i[12];
   assign pp13_o[13] = muler_i[13] & mulcand_i[13];
   assign pp14_o[13] = muler_i[13] & mulcand_i[14];
   assign pp15_o[13] = muler_i[13] & mulcand_i[15];
   assign pp16_o[13] = muler_i[13] & mulcand_i[16];
   assign pp17_o[13] = muler_i[13] & mulcand_i[17];
   assign pp18_o[13] = muler_i[13] & mulcand_i[18];
   assign pp19_o[13] = muler_i[13] & mulcand_i[19];
   assign pp20_o[13] = muler_i[13] & mulcand_i[20];
   assign pp21_o[13] = muler_i[13] & mulcand_i[21];
   assign pp22_o[13] = muler_i[13] & mulcand_i[22];
   assign pp23_o[13] = muler_i[13] & mulcand_i[23];
   assign pp24_o[13] = muler_i[13] & mulcand_i[24];
   assign pp25_o[13] = muler_i[13] & mulcand_i[25];
   assign pp26_o[13] = muler_i[13] & mulcand_i[26];
   assign pp27_o[13] = muler_i[13] & mulcand_i[27];
   assign pp28_o[13] = muler_i[13] & mulcand_i[28];
   assign pp29_o[13] = muler_i[13] & mulcand_i[29];
   assign pp30_o[13] = muler_i[13] & mulcand_i[30];
   assign pp31_o[13] = muler_i[13] & mulcand_i[31];

   assign pp0_o[14]  = muler_i[14] & mulcand_i[0];
   assign pp1_o[14]  = muler_i[14] & mulcand_i[1];
   assign pp2_o[14]  = muler_i[14] & mulcand_i[2];
   assign pp3_o[14]  = muler_i[14] & mulcand_i[3];
   assign pp4_o[14]  = muler_i[14] & mulcand_i[4];
   assign pp5_o[14]  = muler_i[14] & mulcand_i[5];
   assign pp6_o[14]  = muler_i[14] & mulcand_i[6];
   assign pp7_o[14]  = muler_i[14] & mulcand_i[7];
   assign pp8_o[14]  = muler_i[14] & mulcand_i[8];
   assign pp9_o[14]  = muler_i[14] & mulcand_i[9];
   assign pp10_o[14] = muler_i[14] & mulcand_i[10];
   assign pp11_o[14] = muler_i[14] & mulcand_i[11];
   assign pp12_o[14] = muler_i[14] & mulcand_i[12];
   assign pp13_o[14] = muler_i[14] & mulcand_i[13];
   assign pp14_o[14] = muler_i[14] & mulcand_i[14];
   assign pp15_o[14] = muler_i[14] & mulcand_i[15];
   assign pp16_o[14] = muler_i[14] & mulcand_i[16];
   assign pp17_o[14] = muler_i[14] & mulcand_i[17];
   assign pp18_o[14] = muler_i[14] & mulcand_i[18];
   assign pp19_o[14] = muler_i[14] & mulcand_i[19];
   assign pp20_o[14] = muler_i[14] & mulcand_i[20];
   assign pp21_o[14] = muler_i[14] & mulcand_i[21];
   assign pp22_o[14] = muler_i[14] & mulcand_i[22];
   assign pp23_o[14] = muler_i[14] & mulcand_i[23];
   assign pp24_o[14] = muler_i[14] & mulcand_i[24];
   assign pp25_o[14] = muler_i[14] & mulcand_i[25];
   assign pp26_o[14] = muler_i[14] & mulcand_i[26];
   assign pp27_o[14] = muler_i[14] & mulcand_i[27];
   assign pp28_o[14] = muler_i[14] & mulcand_i[28];
   assign pp29_o[14] = muler_i[14] & mulcand_i[29];
   assign pp30_o[14] = muler_i[14] & mulcand_i[30];
   assign pp31_o[14] = muler_i[14] & mulcand_i[31];

   assign pp0_o[15]  = muler_i[15] & mulcand_i[0];
   assign pp1_o[15]  = muler_i[15] & mulcand_i[1];
   assign pp2_o[15]  = muler_i[15] & mulcand_i[2];
   assign pp3_o[15]  = muler_i[15] & mulcand_i[3];
   assign pp4_o[15]  = muler_i[15] & mulcand_i[4];
   assign pp5_o[15]  = muler_i[15] & mulcand_i[5];
   assign pp6_o[15]  = muler_i[15] & mulcand_i[6];
   assign pp7_o[15]  = muler_i[15] & mulcand_i[7];
   assign pp8_o[15]  = muler_i[15] & mulcand_i[8];
   assign pp9_o[15]  = muler_i[15] & mulcand_i[9];
   assign pp10_o[15] = muler_i[15] & mulcand_i[10];
   assign pp11_o[15] = muler_i[15] & mulcand_i[11];
   assign pp12_o[15] = muler_i[15] & mulcand_i[12];
   assign pp13_o[15] = muler_i[15] & mulcand_i[13];
   assign pp14_o[15] = muler_i[15] & mulcand_i[14];
   assign pp15_o[15] = muler_i[15] & mulcand_i[15];
   assign pp16_o[15] = muler_i[15] & mulcand_i[16];
   assign pp17_o[15] = muler_i[15] & mulcand_i[17];
   assign pp18_o[15] = muler_i[15] & mulcand_i[18];
   assign pp19_o[15] = muler_i[15] & mulcand_i[19];
   assign pp20_o[15] = muler_i[15] & mulcand_i[20];
   assign pp21_o[15] = muler_i[15] & mulcand_i[21];
   assign pp22_o[15] = muler_i[15] & mulcand_i[22];
   assign pp23_o[15] = muler_i[15] & mulcand_i[23];
   assign pp24_o[15] = muler_i[15] & mulcand_i[24];
   assign pp25_o[15] = muler_i[15] & mulcand_i[25];
   assign pp26_o[15] = muler_i[15] & mulcand_i[26];
   assign pp27_o[15] = muler_i[15] & mulcand_i[27];
   assign pp28_o[15] = muler_i[15] & mulcand_i[28];
   assign pp29_o[15] = muler_i[15] & mulcand_i[29];
   assign pp30_o[15] = muler_i[15] & mulcand_i[30];
   assign pp31_o[15] = muler_i[15] & mulcand_i[31];

   assign pp0_o[16]  = muler_i[16] & mulcand_i[0];
   assign pp1_o[16]  = muler_i[16] & mulcand_i[1];
   assign pp2_o[16]  = muler_i[16] & mulcand_i[2];
   assign pp3_o[16]  = muler_i[16] & mulcand_i[3];
   assign pp4_o[16]  = muler_i[16] & mulcand_i[4];
   assign pp5_o[16]  = muler_i[16] & mulcand_i[5];
   assign pp6_o[16]  = muler_i[16] & mulcand_i[6];
   assign pp7_o[16]  = muler_i[16] & mulcand_i[7];
   assign pp8_o[16]  = muler_i[16] & mulcand_i[8];
   assign pp9_o[16]  = muler_i[16] & mulcand_i[9];
   assign pp10_o[16] = muler_i[16] & mulcand_i[10];
   assign pp11_o[16] = muler_i[16] & mulcand_i[11];
   assign pp12_o[16] = muler_i[16] & mulcand_i[12];
   assign pp13_o[16] = muler_i[16] & mulcand_i[13];
   assign pp14_o[16] = muler_i[16] & mulcand_i[14];
   assign pp15_o[16] = muler_i[16] & mulcand_i[15];
   assign pp16_o[16] = muler_i[16] & mulcand_i[16];
   assign pp17_o[16] = muler_i[16] & mulcand_i[17];
   assign pp18_o[16] = muler_i[16] & mulcand_i[18];
   assign pp19_o[16] = muler_i[16] & mulcand_i[19];
   assign pp20_o[16] = muler_i[16] & mulcand_i[20];
   assign pp21_o[16] = muler_i[16] & mulcand_i[21];
   assign pp22_o[16] = muler_i[16] & mulcand_i[22];
   assign pp23_o[16] = muler_i[16] & mulcand_i[23];
   assign pp24_o[16] = muler_i[16] & mulcand_i[24];
   assign pp25_o[16] = muler_i[16] & mulcand_i[25];
   assign pp26_o[16] = muler_i[16] & mulcand_i[26];
   assign pp27_o[16] = muler_i[16] & mulcand_i[27];
   assign pp28_o[16] = muler_i[16] & mulcand_i[28];
   assign pp29_o[16] = muler_i[16] & mulcand_i[29];
   assign pp30_o[16] = muler_i[16] & mulcand_i[30];
   assign pp31_o[16] = muler_i[16] & mulcand_i[31];

   assign pp0_o[17]  = muler_i[17] & mulcand_i[0];
   assign pp1_o[17]  = muler_i[17] & mulcand_i[1];
   assign pp2_o[17]  = muler_i[17] & mulcand_i[2];
   assign pp3_o[17]  = muler_i[17] & mulcand_i[3];
   assign pp4_o[17]  = muler_i[17] & mulcand_i[4];
   assign pp5_o[17]  = muler_i[17] & mulcand_i[5];
   assign pp6_o[17]  = muler_i[17] & mulcand_i[6];
   assign pp7_o[17]  = muler_i[17] & mulcand_i[7];
   assign pp8_o[17]  = muler_i[17] & mulcand_i[8];
   assign pp9_o[17]  = muler_i[17] & mulcand_i[9];
   assign pp10_o[17] = muler_i[17] & mulcand_i[10];
   assign pp11_o[17] = muler_i[17] & mulcand_i[11];
   assign pp12_o[17] = muler_i[17] & mulcand_i[12];
   assign pp13_o[17] = muler_i[17] & mulcand_i[13];
   assign pp14_o[17] = muler_i[17] & mulcand_i[14];
   assign pp15_o[17] = muler_i[17] & mulcand_i[15];
   assign pp16_o[17] = muler_i[17] & mulcand_i[16];
   assign pp17_o[17] = muler_i[17] & mulcand_i[17];
   assign pp18_o[17] = muler_i[17] & mulcand_i[18];
   assign pp19_o[17] = muler_i[17] & mulcand_i[19];
   assign pp20_o[17] = muler_i[17] & mulcand_i[20];
   assign pp21_o[17] = muler_i[17] & mulcand_i[21];
   assign pp22_o[17] = muler_i[17] & mulcand_i[22];
   assign pp23_o[17] = muler_i[17] & mulcand_i[23];
   assign pp24_o[17] = muler_i[17] & mulcand_i[24];
   assign pp25_o[17] = muler_i[17] & mulcand_i[25];
   assign pp26_o[17] = muler_i[17] & mulcand_i[26];
   assign pp27_o[17] = muler_i[17] & mulcand_i[27];
   assign pp28_o[17] = muler_i[17] & mulcand_i[28];
   assign pp29_o[17] = muler_i[17] & mulcand_i[29];
   assign pp30_o[17] = muler_i[17] & mulcand_i[30];
   assign pp31_o[17] = muler_i[17] & mulcand_i[31];

   assign pp0_o[18]  = muler_i[18] & mulcand_i[0];
   assign pp1_o[18]  = muler_i[18] & mulcand_i[1];
   assign pp2_o[18]  = muler_i[18] & mulcand_i[2];
   assign pp3_o[18]  = muler_i[18] & mulcand_i[3];
   assign pp4_o[18]  = muler_i[18] & mulcand_i[4];
   assign pp5_o[18]  = muler_i[18] & mulcand_i[5];
   assign pp6_o[18]  = muler_i[18] & mulcand_i[6];
   assign pp7_o[18]  = muler_i[18] & mulcand_i[7];
   assign pp8_o[18]  = muler_i[18] & mulcand_i[8];
   assign pp9_o[18]  = muler_i[18] & mulcand_i[9];
   assign pp10_o[18] = muler_i[18] & mulcand_i[10];
   assign pp11_o[18] = muler_i[18] & mulcand_i[11];
   assign pp12_o[18] = muler_i[18] & mulcand_i[12];
   assign pp13_o[18] = muler_i[18] & mulcand_i[13];
   assign pp14_o[18] = muler_i[18] & mulcand_i[14];
   assign pp15_o[18] = muler_i[18] & mulcand_i[15];
   assign pp16_o[18] = muler_i[18] & mulcand_i[16];
   assign pp17_o[18] = muler_i[18] & mulcand_i[17];
   assign pp18_o[18] = muler_i[18] & mulcand_i[18];
   assign pp19_o[18] = muler_i[18] & mulcand_i[19];
   assign pp20_o[18] = muler_i[18] & mulcand_i[20];
   assign pp21_o[18] = muler_i[18] & mulcand_i[21];
   assign pp22_o[18] = muler_i[18] & mulcand_i[22];
   assign pp23_o[18] = muler_i[18] & mulcand_i[23];
   assign pp24_o[18] = muler_i[18] & mulcand_i[24];
   assign pp25_o[18] = muler_i[18] & mulcand_i[25];
   assign pp26_o[18] = muler_i[18] & mulcand_i[26];
   assign pp27_o[18] = muler_i[18] & mulcand_i[27];
   assign pp28_o[18] = muler_i[18] & mulcand_i[28];
   assign pp29_o[18] = muler_i[18] & mulcand_i[29];
   assign pp30_o[18] = muler_i[18] & mulcand_i[30];
   assign pp31_o[18] = muler_i[18] & mulcand_i[31];

   assign pp0_o[19]  = muler_i[19] & mulcand_i[0];
   assign pp1_o[19]  = muler_i[19] & mulcand_i[1];
   assign pp2_o[19]  = muler_i[19] & mulcand_i[2];
   assign pp3_o[19]  = muler_i[19] & mulcand_i[3];
   assign pp4_o[19]  = muler_i[19] & mulcand_i[4];
   assign pp5_o[19]  = muler_i[19] & mulcand_i[5];
   assign pp6_o[19]  = muler_i[19] & mulcand_i[6];
   assign pp7_o[19]  = muler_i[19] & mulcand_i[7];
   assign pp8_o[19]  = muler_i[19] & mulcand_i[8];
   assign pp9_o[19]  = muler_i[19] & mulcand_i[9];
   assign pp10_o[19] = muler_i[19] & mulcand_i[10];
   assign pp11_o[19] = muler_i[19] & mulcand_i[11];
   assign pp12_o[19] = muler_i[19] & mulcand_i[12];
   assign pp13_o[19] = muler_i[19] & mulcand_i[13];
   assign pp14_o[19] = muler_i[19] & mulcand_i[14];
   assign pp15_o[19] = muler_i[19] & mulcand_i[15];
   assign pp16_o[19] = muler_i[19] & mulcand_i[16];
   assign pp17_o[19] = muler_i[19] & mulcand_i[17];
   assign pp18_o[19] = muler_i[19] & mulcand_i[18];
   assign pp19_o[19] = muler_i[19] & mulcand_i[19];
   assign pp20_o[19] = muler_i[19] & mulcand_i[20];
   assign pp21_o[19] = muler_i[19] & mulcand_i[21];
   assign pp22_o[19] = muler_i[19] & mulcand_i[22];
   assign pp23_o[19] = muler_i[19] & mulcand_i[23];
   assign pp24_o[19] = muler_i[19] & mulcand_i[24];
   assign pp25_o[19] = muler_i[19] & mulcand_i[25];
   assign pp26_o[19] = muler_i[19] & mulcand_i[26];
   assign pp27_o[19] = muler_i[19] & mulcand_i[27];
   assign pp28_o[19] = muler_i[19] & mulcand_i[28];
   assign pp29_o[19] = muler_i[19] & mulcand_i[29];
   assign pp30_o[19] = muler_i[19] & mulcand_i[30];
   assign pp31_o[19] = muler_i[19] & mulcand_i[31];

   assign pp0_o[20]  = muler_i[20] & mulcand_i[0];
   assign pp1_o[20]  = muler_i[20] & mulcand_i[1];
   assign pp2_o[20]  = muler_i[20] & mulcand_i[2];
   assign pp3_o[20]  = muler_i[20] & mulcand_i[3];
   assign pp4_o[20]  = muler_i[20] & mulcand_i[4];
   assign pp5_o[20]  = muler_i[20] & mulcand_i[5];
   assign pp6_o[20]  = muler_i[20] & mulcand_i[6];
   assign pp7_o[20]  = muler_i[20] & mulcand_i[7];
   assign pp8_o[20]  = muler_i[20] & mulcand_i[8];
   assign pp9_o[20]  = muler_i[20] & mulcand_i[9];
   assign pp10_o[20] = muler_i[20] & mulcand_i[10];
   assign pp11_o[20] = muler_i[20] & mulcand_i[11];
   assign pp12_o[20] = muler_i[20] & mulcand_i[12];
   assign pp13_o[20] = muler_i[20] & mulcand_i[13];
   assign pp14_o[20] = muler_i[20] & mulcand_i[14];
   assign pp15_o[20] = muler_i[20] & mulcand_i[15];
   assign pp16_o[20] = muler_i[20] & mulcand_i[16];
   assign pp17_o[20] = muler_i[20] & mulcand_i[17];
   assign pp18_o[20] = muler_i[20] & mulcand_i[18];
   assign pp19_o[20] = muler_i[20] & mulcand_i[19];
   assign pp20_o[20] = muler_i[20] & mulcand_i[20];
   assign pp21_o[20] = muler_i[20] & mulcand_i[21];
   assign pp22_o[20] = muler_i[20] & mulcand_i[22];
   assign pp23_o[20] = muler_i[20] & mulcand_i[23];
   assign pp24_o[20] = muler_i[20] & mulcand_i[24];
   assign pp25_o[20] = muler_i[20] & mulcand_i[25];
   assign pp26_o[20] = muler_i[20] & mulcand_i[26];
   assign pp27_o[20] = muler_i[20] & mulcand_i[27];
   assign pp28_o[20] = muler_i[20] & mulcand_i[28];
   assign pp29_o[20] = muler_i[20] & mulcand_i[29];
   assign pp30_o[20] = muler_i[20] & mulcand_i[30];
   assign pp31_o[20] = muler_i[20] & mulcand_i[31];

   assign pp0_o[21]  = muler_i[21] & mulcand_i[0];
   assign pp1_o[21]  = muler_i[21] & mulcand_i[1];
   assign pp2_o[21]  = muler_i[21] & mulcand_i[2];
   assign pp3_o[21]  = muler_i[21] & mulcand_i[3];
   assign pp4_o[21]  = muler_i[21] & mulcand_i[4];
   assign pp5_o[21]  = muler_i[21] & mulcand_i[5];
   assign pp6_o[21]  = muler_i[21] & mulcand_i[6];
   assign pp7_o[21]  = muler_i[21] & mulcand_i[7];
   assign pp8_o[21]  = muler_i[21] & mulcand_i[8];
   assign pp9_o[21]  = muler_i[21] & mulcand_i[9];
   assign pp10_o[21] = muler_i[21] & mulcand_i[10];
   assign pp11_o[21] = muler_i[21] & mulcand_i[11];
   assign pp12_o[21] = muler_i[21] & mulcand_i[12];
   assign pp13_o[21] = muler_i[21] & mulcand_i[13];
   assign pp14_o[21] = muler_i[21] & mulcand_i[14];
   assign pp15_o[21] = muler_i[21] & mulcand_i[15];
   assign pp16_o[21] = muler_i[21] & mulcand_i[16];
   assign pp17_o[21] = muler_i[21] & mulcand_i[17];
   assign pp18_o[21] = muler_i[21] & mulcand_i[18];
   assign pp19_o[21] = muler_i[21] & mulcand_i[19];
   assign pp20_o[21] = muler_i[21] & mulcand_i[20];
   assign pp21_o[21] = muler_i[21] & mulcand_i[21];
   assign pp22_o[21] = muler_i[21] & mulcand_i[22];
   assign pp23_o[21] = muler_i[21] & mulcand_i[23];
   assign pp24_o[21] = muler_i[21] & mulcand_i[24];
   assign pp25_o[21] = muler_i[21] & mulcand_i[25];
   assign pp26_o[21] = muler_i[21] & mulcand_i[26];
   assign pp27_o[21] = muler_i[21] & mulcand_i[27];
   assign pp28_o[21] = muler_i[21] & mulcand_i[28];
   assign pp29_o[21] = muler_i[21] & mulcand_i[29];
   assign pp30_o[21] = muler_i[21] & mulcand_i[30];
   assign pp31_o[21] = muler_i[21] & mulcand_i[31];
      
   assign pp0_o[22]  = muler_i[22] & mulcand_i[0];
   assign pp1_o[22]  = muler_i[22] & mulcand_i[1];
   assign pp2_o[22]  = muler_i[22] & mulcand_i[2];
   assign pp3_o[22]  = muler_i[22] & mulcand_i[3];
   assign pp4_o[22]  = muler_i[22] & mulcand_i[4];
   assign pp5_o[22]  = muler_i[22] & mulcand_i[5];
   assign pp6_o[22]  = muler_i[22] & mulcand_i[6];
   assign pp7_o[22]  = muler_i[22] & mulcand_i[7];
   assign pp8_o[22]  = muler_i[22] & mulcand_i[8];
   assign pp9_o[22]  = muler_i[22] & mulcand_i[9];
   assign pp10_o[22] = muler_i[22] & mulcand_i[10];
   assign pp11_o[22] = muler_i[22] & mulcand_i[11];
   assign pp12_o[22] = muler_i[22] & mulcand_i[12];
   assign pp13_o[22] = muler_i[22] & mulcand_i[13];
   assign pp14_o[22] = muler_i[22] & mulcand_i[14];
   assign pp15_o[22] = muler_i[22] & mulcand_i[15];
   assign pp16_o[22] = muler_i[22] & mulcand_i[16];
   assign pp17_o[22] = muler_i[22] & mulcand_i[17];
   assign pp18_o[22] = muler_i[22] & mulcand_i[18];
   assign pp19_o[22] = muler_i[22] & mulcand_i[19];
   assign pp20_o[22] = muler_i[22] & mulcand_i[20];
   assign pp21_o[22] = muler_i[22] & mulcand_i[21];
   assign pp22_o[22] = muler_i[22] & mulcand_i[22];
   assign pp23_o[22] = muler_i[22] & mulcand_i[23];
   assign pp24_o[22] = muler_i[22] & mulcand_i[24];
   assign pp25_o[22] = muler_i[22] & mulcand_i[25];
   assign pp26_o[22] = muler_i[22] & mulcand_i[26];
   assign pp27_o[22] = muler_i[22] & mulcand_i[27];
   assign pp28_o[22] = muler_i[22] & mulcand_i[28];
   assign pp29_o[22] = muler_i[22] & mulcand_i[29];
   assign pp30_o[22] = muler_i[22] & mulcand_i[30];
   assign pp31_o[22] = muler_i[22] & mulcand_i[31];

   assign pp0_o[23]  = muler_i[23] & mulcand_i[0];
   assign pp1_o[23]  = muler_i[23] & mulcand_i[1];
   assign pp2_o[23]  = muler_i[23] & mulcand_i[2];
   assign pp3_o[23]  = muler_i[23] & mulcand_i[3];
   assign pp4_o[23]  = muler_i[23] & mulcand_i[4];
   assign pp5_o[23]  = muler_i[23] & mulcand_i[5];
   assign pp6_o[23]  = muler_i[23] & mulcand_i[6];
   assign pp7_o[23]  = muler_i[23] & mulcand_i[7];
   assign pp8_o[23]  = muler_i[23] & mulcand_i[8];
   assign pp9_o[23]  = muler_i[23] & mulcand_i[9];
   assign pp10_o[23] = muler_i[23] & mulcand_i[10];
   assign pp11_o[23] = muler_i[23] & mulcand_i[11];
   assign pp12_o[23] = muler_i[23] & mulcand_i[12];
   assign pp13_o[23] = muler_i[23] & mulcand_i[13];
   assign pp14_o[23] = muler_i[23] & mulcand_i[14];
   assign pp15_o[23] = muler_i[23] & mulcand_i[15];
   assign pp16_o[23] = muler_i[23] & mulcand_i[16];
   assign pp17_o[23] = muler_i[23] & mulcand_i[17];
   assign pp18_o[23] = muler_i[23] & mulcand_i[18];
   assign pp19_o[23] = muler_i[23] & mulcand_i[19];
   assign pp20_o[23] = muler_i[23] & mulcand_i[20];
   assign pp21_o[23] = muler_i[23] & mulcand_i[21];
   assign pp22_o[23] = muler_i[23] & mulcand_i[22];
   assign pp23_o[23] = muler_i[23] & mulcand_i[23];
   assign pp24_o[23] = muler_i[23] & mulcand_i[24];
   assign pp25_o[23] = muler_i[23] & mulcand_i[25];
   assign pp26_o[23] = muler_i[23] & mulcand_i[26];
   assign pp27_o[23] = muler_i[23] & mulcand_i[27];
   assign pp28_o[23] = muler_i[23] & mulcand_i[28];
   assign pp29_o[23] = muler_i[23] & mulcand_i[29];
   assign pp30_o[23] = muler_i[23] & mulcand_i[30];
   assign pp31_o[23] = muler_i[23] & mulcand_i[31];

   assign pp0_o[24]  = muler_i[24] & mulcand_i[0];
   assign pp1_o[24]  = muler_i[24] & mulcand_i[1];
   assign pp2_o[24]  = muler_i[24] & mulcand_i[2];
   assign pp3_o[24]  = muler_i[24] & mulcand_i[3];
   assign pp4_o[24]  = muler_i[24] & mulcand_i[4];
   assign pp5_o[24]  = muler_i[24] & mulcand_i[5];
   assign pp6_o[24]  = muler_i[24] & mulcand_i[6];
   assign pp7_o[24]  = muler_i[24] & mulcand_i[7];
   assign pp8_o[24]  = muler_i[24] & mulcand_i[8];
   assign pp9_o[24]  = muler_i[24] & mulcand_i[9];
   assign pp10_o[24] = muler_i[24] & mulcand_i[10];
   assign pp11_o[24] = muler_i[24] & mulcand_i[11];
   assign pp12_o[24] = muler_i[24] & mulcand_i[12];
   assign pp13_o[24] = muler_i[24] & mulcand_i[13];
   assign pp14_o[24] = muler_i[24] & mulcand_i[14];
   assign pp15_o[24] = muler_i[24] & mulcand_i[15];
   assign pp16_o[24] = muler_i[24] & mulcand_i[16];
   assign pp17_o[24] = muler_i[24] & mulcand_i[17];
   assign pp18_o[24] = muler_i[24] & mulcand_i[18];
   assign pp19_o[24] = muler_i[24] & mulcand_i[19];
   assign pp20_o[24] = muler_i[24] & mulcand_i[20];
   assign pp21_o[24] = muler_i[24] & mulcand_i[21];
   assign pp22_o[24] = muler_i[24] & mulcand_i[22];
   assign pp23_o[24] = muler_i[24] & mulcand_i[23];
   assign pp24_o[24] = muler_i[24] & mulcand_i[24];
   assign pp25_o[24] = muler_i[24] & mulcand_i[25];
   assign pp26_o[24] = muler_i[24] & mulcand_i[26];
   assign pp27_o[24] = muler_i[24] & mulcand_i[27];
   assign pp28_o[24] = muler_i[24] & mulcand_i[28];
   assign pp29_o[24] = muler_i[24] & mulcand_i[29];
   assign pp30_o[24] = muler_i[24] & mulcand_i[30];
   assign pp31_o[24] = muler_i[24] & mulcand_i[31];

   assign pp0_o[25]  = muler_i[25] & mulcand_i[0];
   assign pp1_o[25]  = muler_i[25] & mulcand_i[1];
   assign pp2_o[25]  = muler_i[25] & mulcand_i[2];
   assign pp3_o[25]  = muler_i[25] & mulcand_i[3];
   assign pp4_o[25]  = muler_i[25] & mulcand_i[4];
   assign pp5_o[25]  = muler_i[25] & mulcand_i[5];
   assign pp6_o[25]  = muler_i[25] & mulcand_i[6];
   assign pp7_o[25]  = muler_i[25] & mulcand_i[7];
   assign pp8_o[25]  = muler_i[25] & mulcand_i[8];
   assign pp9_o[25]  = muler_i[25] & mulcand_i[9];
   assign pp10_o[25] = muler_i[25] & mulcand_i[10];
   assign pp11_o[25] = muler_i[25] & mulcand_i[11];
   assign pp12_o[25] = muler_i[25] & mulcand_i[12];
   assign pp13_o[25] = muler_i[25] & mulcand_i[13];
   assign pp14_o[25] = muler_i[25] & mulcand_i[14];
   assign pp15_o[25] = muler_i[25] & mulcand_i[15];
   assign pp16_o[25] = muler_i[25] & mulcand_i[16];
   assign pp17_o[25] = muler_i[25] & mulcand_i[17];
   assign pp18_o[25] = muler_i[25] & mulcand_i[18];
   assign pp19_o[25] = muler_i[25] & mulcand_i[19];
   assign pp20_o[25] = muler_i[25] & mulcand_i[20];
   assign pp21_o[25] = muler_i[25] & mulcand_i[21];
   assign pp22_o[25] = muler_i[25] & mulcand_i[22];
   assign pp23_o[25] = muler_i[25] & mulcand_i[23];
   assign pp24_o[25] = muler_i[25] & mulcand_i[24];
   assign pp25_o[25] = muler_i[25] & mulcand_i[25];
   assign pp26_o[25] = muler_i[25] & mulcand_i[26];
   assign pp27_o[25] = muler_i[25] & mulcand_i[27];
   assign pp28_o[25] = muler_i[25] & mulcand_i[28];
   assign pp29_o[25] = muler_i[25] & mulcand_i[29];
   assign pp30_o[25] = muler_i[25] & mulcand_i[30];
   assign pp31_o[25] = muler_i[25] & mulcand_i[31];

   assign pp0_o[26]  = muler_i[26] & mulcand_i[0];
   assign pp1_o[26]  = muler_i[26] & mulcand_i[1];
   assign pp2_o[26]  = muler_i[26] & mulcand_i[2];
   assign pp3_o[26]  = muler_i[26] & mulcand_i[3];
   assign pp4_o[26]  = muler_i[26] & mulcand_i[4];
   assign pp5_o[26]  = muler_i[26] & mulcand_i[5];
   assign pp6_o[26]  = muler_i[26] & mulcand_i[6];
   assign pp7_o[26]  = muler_i[26] & mulcand_i[7];
   assign pp8_o[26]  = muler_i[26] & mulcand_i[8];
   assign pp9_o[26]  = muler_i[26] & mulcand_i[9];
   assign pp10_o[26] = muler_i[26] & mulcand_i[10];
   assign pp11_o[26] = muler_i[26] & mulcand_i[11];
   assign pp12_o[26] = muler_i[26] & mulcand_i[12];
   assign pp13_o[26] = muler_i[26] & mulcand_i[13];
   assign pp14_o[26] = muler_i[26] & mulcand_i[14];
   assign pp15_o[26] = muler_i[26] & mulcand_i[15];
   assign pp16_o[26] = muler_i[26] & mulcand_i[16];
   assign pp17_o[26] = muler_i[26] & mulcand_i[17];
   assign pp18_o[26] = muler_i[26] & mulcand_i[18];
   assign pp19_o[26] = muler_i[26] & mulcand_i[19];
   assign pp20_o[26] = muler_i[26] & mulcand_i[20];
   assign pp21_o[26] = muler_i[26] & mulcand_i[21];
   assign pp22_o[26] = muler_i[26] & mulcand_i[22];
   assign pp23_o[26] = muler_i[26] & mulcand_i[23];
   assign pp24_o[26] = muler_i[26] & mulcand_i[24];
   assign pp25_o[26] = muler_i[26] & mulcand_i[25];
   assign pp26_o[26] = muler_i[26] & mulcand_i[26];
   assign pp27_o[26] = muler_i[26] & mulcand_i[27];
   assign pp28_o[26] = muler_i[26] & mulcand_i[28];
   assign pp29_o[26] = muler_i[26] & mulcand_i[29];
   assign pp30_o[26] = muler_i[26] & mulcand_i[30];
   assign pp31_o[26] = muler_i[26] & mulcand_i[31];

   assign pp0_o[27]  = muler_i[27] & mulcand_i[0];
   assign pp1_o[27]  = muler_i[27] & mulcand_i[1];
   assign pp2_o[27]  = muler_i[27] & mulcand_i[2];
   assign pp3_o[27]  = muler_i[27] & mulcand_i[3];
   assign pp4_o[27]  = muler_i[27] & mulcand_i[4];
   assign pp5_o[27]  = muler_i[27] & mulcand_i[5];
   assign pp6_o[27]  = muler_i[27] & mulcand_i[6];
   assign pp7_o[27]  = muler_i[27] & mulcand_i[7];
   assign pp8_o[27]  = muler_i[27] & mulcand_i[8];
   assign pp9_o[27]  = muler_i[27] & mulcand_i[9];
   assign pp10_o[27] = muler_i[27] & mulcand_i[10];
   assign pp11_o[27] = muler_i[27] & mulcand_i[11];
   assign pp12_o[27] = muler_i[27] & mulcand_i[12];
   assign pp13_o[27] = muler_i[27] & mulcand_i[13];
   assign pp14_o[27] = muler_i[27] & mulcand_i[14];
   assign pp15_o[27] = muler_i[27] & mulcand_i[15];
   assign pp16_o[27] = muler_i[27] & mulcand_i[16];
   assign pp17_o[27] = muler_i[27] & mulcand_i[17];
   assign pp18_o[27] = muler_i[27] & mulcand_i[18];
   assign pp19_o[27] = muler_i[27] & mulcand_i[19];
   assign pp20_o[27] = muler_i[27] & mulcand_i[20];
   assign pp21_o[27] = muler_i[27] & mulcand_i[21];
   assign pp22_o[27] = muler_i[27] & mulcand_i[22];
   assign pp23_o[27] = muler_i[27] & mulcand_i[23];
   assign pp24_o[27] = muler_i[27] & mulcand_i[24];
   assign pp25_o[27] = muler_i[27] & mulcand_i[25];
   assign pp26_o[27] = muler_i[27] & mulcand_i[26];
   assign pp27_o[27] = muler_i[27] & mulcand_i[27];
   assign pp28_o[27] = muler_i[27] & mulcand_i[28];
   assign pp29_o[27] = muler_i[27] & mulcand_i[29];
   assign pp30_o[27] = muler_i[27] & mulcand_i[30];
   assign pp31_o[27] = muler_i[27] & mulcand_i[31];

   assign pp0_o[28]  = muler_i[28] & mulcand_i[0];
   assign pp1_o[28]  = muler_i[28] & mulcand_i[1];
   assign pp2_o[28]  = muler_i[28] & mulcand_i[2];
   assign pp3_o[28]  = muler_i[28] & mulcand_i[3];
   assign pp4_o[28]  = muler_i[28] & mulcand_i[4];
   assign pp5_o[28]  = muler_i[28] & mulcand_i[5];
   assign pp6_o[28]  = muler_i[28] & mulcand_i[6];
   assign pp7_o[28]  = muler_i[28] & mulcand_i[7];
   assign pp8_o[28]  = muler_i[28] & mulcand_i[8];
   assign pp9_o[28]  = muler_i[28] & mulcand_i[9];
   assign pp10_o[28] = muler_i[28] & mulcand_i[10];
   assign pp11_o[28] = muler_i[28] & mulcand_i[11];
   assign pp12_o[28] = muler_i[28] & mulcand_i[12];
   assign pp13_o[28] = muler_i[28] & mulcand_i[13];
   assign pp14_o[28] = muler_i[28] & mulcand_i[14];
   assign pp15_o[28] = muler_i[28] & mulcand_i[15];
   assign pp16_o[28] = muler_i[28] & mulcand_i[16];
   assign pp17_o[28] = muler_i[28] & mulcand_i[17];
   assign pp18_o[28] = muler_i[28] & mulcand_i[18];
   assign pp19_o[28] = muler_i[28] & mulcand_i[19];
   assign pp20_o[28] = muler_i[28] & mulcand_i[20];
   assign pp21_o[28] = muler_i[28] & mulcand_i[21];
   assign pp22_o[28] = muler_i[28] & mulcand_i[22];
   assign pp23_o[28] = muler_i[28] & mulcand_i[23];
   assign pp24_o[28] = muler_i[28] & mulcand_i[24];
   assign pp25_o[28] = muler_i[28] & mulcand_i[25];
   assign pp26_o[28] = muler_i[28] & mulcand_i[26];
   assign pp27_o[28] = muler_i[28] & mulcand_i[27];
   assign pp28_o[28] = muler_i[28] & mulcand_i[28];
   assign pp29_o[28] = muler_i[28] & mulcand_i[29];
   assign pp30_o[28] = muler_i[28] & mulcand_i[30];
   assign pp31_o[28] = muler_i[28] & mulcand_i[31];

   assign pp0_o[29]  = muler_i[29] & mulcand_i[0];
   assign pp1_o[29]  = muler_i[29] & mulcand_i[1];
   assign pp2_o[29]  = muler_i[29] & mulcand_i[2];
   assign pp3_o[29]  = muler_i[29] & mulcand_i[3];
   assign pp4_o[29]  = muler_i[29] & mulcand_i[4];
   assign pp5_o[29]  = muler_i[29] & mulcand_i[5];
   assign pp6_o[29]  = muler_i[29] & mulcand_i[6];
   assign pp7_o[29]  = muler_i[29] & mulcand_i[7];
   assign pp8_o[29]  = muler_i[29] & mulcand_i[8];
   assign pp9_o[29]  = muler_i[29] & mulcand_i[9];
   assign pp10_o[29] = muler_i[29] & mulcand_i[10];
   assign pp11_o[29] = muler_i[29] & mulcand_i[11];
   assign pp12_o[29] = muler_i[29] & mulcand_i[12];
   assign pp13_o[29] = muler_i[29] & mulcand_i[13];
   assign pp14_o[29] = muler_i[29] & mulcand_i[14];
   assign pp15_o[29] = muler_i[29] & mulcand_i[15];
   assign pp16_o[29] = muler_i[29] & mulcand_i[16];
   assign pp17_o[29] = muler_i[29] & mulcand_i[17];
   assign pp18_o[29] = muler_i[29] & mulcand_i[18];
   assign pp19_o[29] = muler_i[29] & mulcand_i[19];
   assign pp20_o[29] = muler_i[29] & mulcand_i[20];
   assign pp21_o[29] = muler_i[29] & mulcand_i[21];
   assign pp22_o[29] = muler_i[29] & mulcand_i[22];
   assign pp23_o[29] = muler_i[29] & mulcand_i[23];
   assign pp24_o[29] = muler_i[29] & mulcand_i[24];
   assign pp25_o[29] = muler_i[29] & mulcand_i[25];
   assign pp26_o[29] = muler_i[29] & mulcand_i[26];
   assign pp27_o[29] = muler_i[29] & mulcand_i[27];
   assign pp28_o[29] = muler_i[29] & mulcand_i[28];
   assign pp29_o[29] = muler_i[29] & mulcand_i[29];
   assign pp30_o[29] = muler_i[29] & mulcand_i[30];
   assign pp31_o[29] = muler_i[29] & mulcand_i[31];

   assign pp0_o[30]  = muler_i[30] & mulcand_i[0];
   assign pp1_o[30]  = muler_i[30] & mulcand_i[1];
   assign pp2_o[30]  = muler_i[30] & mulcand_i[2];
   assign pp3_o[30]  = muler_i[30] & mulcand_i[3];
   assign pp4_o[30]  = muler_i[30] & mulcand_i[4];
   assign pp5_o[30]  = muler_i[30] & mulcand_i[5];
   assign pp6_o[30]  = muler_i[30] & mulcand_i[6];
   assign pp7_o[30]  = muler_i[30] & mulcand_i[7];
   assign pp8_o[30]  = muler_i[30] & mulcand_i[8];
   assign pp9_o[30]  = muler_i[30] & mulcand_i[9];
   assign pp10_o[30] = muler_i[30] & mulcand_i[10];
   assign pp11_o[30] = muler_i[30] & mulcand_i[11];
   assign pp12_o[30] = muler_i[30] & mulcand_i[12];
   assign pp13_o[30] = muler_i[30] & mulcand_i[13];
   assign pp14_o[30] = muler_i[30] & mulcand_i[14];
   assign pp15_o[30] = muler_i[30] & mulcand_i[15];
   assign pp16_o[30] = muler_i[30] & mulcand_i[16];
   assign pp17_o[30] = muler_i[30] & mulcand_i[17];
   assign pp18_o[30] = muler_i[30] & mulcand_i[18];
   assign pp19_o[30] = muler_i[30] & mulcand_i[19];
   assign pp20_o[30] = muler_i[30] & mulcand_i[20];
   assign pp21_o[30] = muler_i[30] & mulcand_i[21];
   assign pp22_o[30] = muler_i[30] & mulcand_i[22];
   assign pp23_o[30] = muler_i[30] & mulcand_i[23];
   assign pp24_o[30] = muler_i[30] & mulcand_i[24];
   assign pp25_o[30] = muler_i[30] & mulcand_i[25];
   assign pp26_o[30] = muler_i[30] & mulcand_i[26];
   assign pp27_o[30] = muler_i[30] & mulcand_i[27];
   assign pp28_o[30] = muler_i[30] & mulcand_i[28];
   assign pp29_o[30] = muler_i[30] & mulcand_i[29];
   assign pp30_o[30] = muler_i[30] & mulcand_i[30];
   assign pp31_o[30] = muler_i[30] & mulcand_i[31];

   assign pp0_o[31]  = muler_i[31] & mulcand_i[0];
   assign pp1_o[31]  = muler_i[31] & mulcand_i[1];
   assign pp2_o[31]  = muler_i[31] & mulcand_i[2];
   assign pp3_o[31]  = muler_i[31] & mulcand_i[3];
   assign pp4_o[31]  = muler_i[31] & mulcand_i[4];
   assign pp5_o[31]  = muler_i[31] & mulcand_i[5];
   assign pp6_o[31]  = muler_i[31] & mulcand_i[6];
   assign pp7_o[31]  = muler_i[31] & mulcand_i[7];
   assign pp8_o[31]  = muler_i[31] & mulcand_i[8];
   assign pp9_o[31]  = muler_i[31] & mulcand_i[9];
   assign pp10_o[31] = muler_i[31] & mulcand_i[10];
   assign pp11_o[31] = muler_i[31] & mulcand_i[11];
   assign pp12_o[31] = muler_i[31] & mulcand_i[12];
   assign pp13_o[31] = muler_i[31] & mulcand_i[13];
   assign pp14_o[31] = muler_i[31] & mulcand_i[14];
   assign pp15_o[31] = muler_i[31] & mulcand_i[15];
   assign pp16_o[31] = muler_i[31] & mulcand_i[16];
   assign pp17_o[31] = muler_i[31] & mulcand_i[17];
   assign pp18_o[31] = muler_i[31] & mulcand_i[18];
   assign pp19_o[31] = muler_i[31] & mulcand_i[19];
   assign pp20_o[31] = muler_i[31] & mulcand_i[20];
   assign pp21_o[31] = muler_i[31] & mulcand_i[21];
   assign pp22_o[31] = muler_i[31] & mulcand_i[22];
   assign pp23_o[31] = muler_i[31] & mulcand_i[23];
   assign pp24_o[31] = muler_i[31] & mulcand_i[24];
   assign pp25_o[31] = muler_i[31] & mulcand_i[25];
   assign pp26_o[31] = muler_i[31] & mulcand_i[26];
   assign pp27_o[31] = muler_i[31] & mulcand_i[27];
   assign pp28_o[31] = muler_i[31] & mulcand_i[28];
   assign pp29_o[31] = muler_i[31] & mulcand_i[29];
   assign pp30_o[31] = muler_i[31] & mulcand_i[30];
   assign pp31_o[31] = muler_i[31] & mulcand_i[31];

endmodule
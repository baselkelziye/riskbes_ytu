
function   mult (input  [3:0] address1, input [3:0] address2);

parameter [7:0] ROM[255:0] = {
		8'd225, 	 // 15 x 15
		8'd210, 	 // 15 x 14
		8'd195, 	 // 15 x 13
		8'd180, 	 // 15 x 12
		8'd165, 	 // 15 x 11
		8'd150, 	 // 15 x 10
		8'd135, 	 // 15 x 9
		8'd120, 	 // 15 x 8
		8'd105, 	 // 15 x 7
		8'd90, 	 // 15 x 6
		8'd75, 	 // 15 x 5
		8'd60, 	 // 15 x 4
		8'd45, 	 // 15 x 3
		8'd30, 	 // 15 x 2
		8'd15, 	 // 15 x 1
		8'd0, 	 // 15 x 0
		8'd210, 	 // 14 x 15
		8'd196, 	 // 14 x 14
		8'd182, 	 // 14 x 13
		8'd168, 	 // 14 x 12
		8'd154, 	 // 14 x 11
		8'd140, 	 // 14 x 10
		8'd126, 	 // 14 x 9
		8'd112, 	 // 14 x 8
		8'd98, 	 // 14 x 7
		8'd84, 	 // 14 x 6
		8'd70, 	 // 14 x 5
		8'd56, 	 // 14 x 4
		8'd42, 	 // 14 x 3
		8'd28, 	 // 14 x 2
		8'd14, 	 // 14 x 1
		8'd0, 	 // 14 x 0
		8'd195, 	 // 13 x 15
		8'd182, 	 // 13 x 14
		8'd169, 	 // 13 x 13
		8'd156, 	 // 13 x 12
		8'd143, 	 // 13 x 11
		8'd130, 	 // 13 x 10
		8'd117, 	 // 13 x 9
		8'd104, 	 // 13 x 8
		8'd91, 	 // 13 x 7
		8'd78, 	 // 13 x 6
		8'd65, 	 // 13 x 5
		8'd52, 	 // 13 x 4
		8'd39, 	 // 13 x 3
		8'd26, 	 // 13 x 2
		8'd13, 	 // 13 x 1
		8'd0, 	 // 13 x 0
		8'd180, 	 // 12 x 15
		8'd168, 	 // 12 x 14
		8'd156, 	 // 12 x 13
		8'd144, 	 // 12 x 12
		8'd132, 	 // 12 x 11
		8'd120, 	 // 12 x 10
		8'd108, 	 // 12 x 9
		8'd96, 	 // 12 x 8
		8'd84, 	 // 12 x 7
		8'd72, 	 // 12 x 6
		8'd60, 	 // 12 x 5
		8'd48, 	 // 12 x 4
		8'd36, 	 // 12 x 3
		8'd24, 	 // 12 x 2
		8'd12, 	 // 12 x 1
		8'd0, 	 // 12 x 0
		8'd165, 	 // 11 x 15
		8'd154, 	 // 11 x 14
		8'd143, 	 // 11 x 13
		8'd132, 	 // 11 x 12
		8'd121, 	 // 11 x 11
		8'd110, 	 // 11 x 10
		8'd99, 	 // 11 x 9
		8'd88, 	 // 11 x 8
		8'd77, 	 // 11 x 7
		8'd66, 	 // 11 x 6
		8'd55, 	 // 11 x 5
		8'd44, 	 // 11 x 4
		8'd33, 	 // 11 x 3
		8'd22, 	 // 11 x 2
		8'd11, 	 // 11 x 1
		8'd0, 	 // 11 x 0
		8'd150, 	 // 10 x 15
		8'd140, 	 // 10 x 14
		8'd130, 	 // 10 x 13
		8'd120, 	 // 10 x 12
		8'd110, 	 // 10 x 11
		8'd100, 	 // 10 x 10
		8'd90, 	 // 10 x 9
		8'd80, 	 // 10 x 8
		8'd70, 	 // 10 x 7
		8'd60, 	 // 10 x 6
		8'd50, 	 // 10 x 5
		8'd40, 	 // 10 x 4
		8'd30, 	 // 10 x 3
		8'd20, 	 // 10 x 2
		8'd10, 	 // 10 x 1
		8'd0, 	 // 10 x 0
		8'd135, 	 // 9 x 15
		8'd126, 	 // 9 x 14
		8'd117, 	 // 9 x 13
		8'd108, 	 // 9 x 12
		8'd99, 	 // 9 x 11
		8'd90, 	 // 9 x 10
		8'd81, 	 // 9 x 9
		8'd72, 	 // 9 x 8
		8'd63, 	 // 9 x 7
		8'd54, 	 // 9 x 6
		8'd45, 	 // 9 x 5
		8'd36, 	 // 9 x 4
		8'd27, 	 // 9 x 3
		8'd18, 	 // 9 x 2
		8'd9, 	 // 9 x 1
		8'd0, 	 // 9 x 0
		8'd120, 	 // 8 x 15
		8'd112, 	 // 8 x 14
		8'd104, 	 // 8 x 13
		8'd96, 	 // 8 x 12
		8'd88, 	 // 8 x 11
		8'd80, 	 // 8 x 10
		8'd72, 	 // 8 x 9
		8'd64, 	 // 8 x 8
		8'd56, 	 // 8 x 7
		8'd48, 	 // 8 x 6
		8'd40, 	 // 8 x 5
		8'd32, 	 // 8 x 4
		8'd24, 	 // 8 x 3
		8'd16, 	 // 8 x 2
		8'd8, 	 // 8 x 1
		8'd0, 	 // 8 x 0
		8'd105, 	 // 7 x 15
		8'd98, 	 // 7 x 14
		8'd91, 	 // 7 x 13
		8'd84, 	 // 7 x 12
		8'd77, 	 // 7 x 11
		8'd70, 	 // 7 x 10
		8'd63, 	 // 7 x 9
		8'd56, 	 // 7 x 8
		8'd49, 	 // 7 x 7
		8'd42, 	 // 7 x 6
		8'd35, 	 // 7 x 5
		8'd28, 	 // 7 x 4
		8'd21, 	 // 7 x 3
		8'd14, 	 // 7 x 2
		8'd7, 	 // 7 x 1
		8'd0, 	 // 7 x 0
		8'd90, 	 // 6 x 15
		8'd84, 	 // 6 x 14
		8'd78, 	 // 6 x 13
		8'd72, 	 // 6 x 12
		8'd66, 	 // 6 x 11
		8'd60, 	 // 6 x 10
		8'd54, 	 // 6 x 9
		8'd48, 	 // 6 x 8
		8'd42, 	 // 6 x 7
		8'd36, 	 // 6 x 6
		8'd30, 	 // 6 x 5
		8'd24, 	 // 6 x 4
		8'd18, 	 // 6 x 3
		8'd12, 	 // 6 x 2
		8'd6, 	 // 6 x 1
		8'd0, 	 // 6 x 0
		8'd75, 	 // 5 x 15
		8'd70, 	 // 5 x 14
		8'd65, 	 // 5 x 13
		8'd60, 	 // 5 x 12
		8'd55, 	 // 5 x 11
		8'd50, 	 // 5 x 10
		8'd45, 	 // 5 x 9
		8'd40, 	 // 5 x 8
		8'd35, 	 // 5 x 7
		8'd30, 	 // 5 x 6
		8'd25, 	 // 5 x 5
		8'd20, 	 // 5 x 4
		8'd15, 	 // 5 x 3
		8'd10, 	 // 5 x 2
		8'd5, 	 // 5 x 1
		8'd0, 	 // 5 x 0
		8'd60, 	 // 4 x 15
		8'd56, 	 // 4 x 14
		8'd52, 	 // 4 x 13
		8'd48, 	 // 4 x 12
		8'd44, 	 // 4 x 11
		8'd40, 	 // 4 x 10
		8'd36, 	 // 4 x 9
		8'd32, 	 // 4 x 8
		8'd28, 	 // 4 x 7
		8'd24, 	 // 4 x 6
		8'd20, 	 // 4 x 5
		8'd16, 	 // 4 x 4
		8'd12, 	 // 4 x 3
		8'd8, 	 // 4 x 2
		8'd4, 	 // 4 x 1
		8'd0, 	 // 4 x 0
		8'd45, 	 // 3 x 15
		8'd42, 	 // 3 x 14
		8'd39, 	 // 3 x 13
		8'd36, 	 // 3 x 12
		8'd33, 	 // 3 x 11
		8'd30, 	 // 3 x 10
		8'd27, 	 // 3 x 9
		8'd24, 	 // 3 x 8
		8'd21, 	 // 3 x 7
		8'd18, 	 // 3 x 6
		8'd15, 	 // 3 x 5
		8'd12, 	 // 3 x 4
		8'd9, 	 // 3 x 3
		8'd6, 	 // 3 x 2
		8'd3, 	 // 3 x 1
		8'd0, 	 // 3 x 0
		8'd30, 	 // 2 x 15
		8'd28, 	 // 2 x 14
		8'd26, 	 // 2 x 13
		8'd24, 	 // 2 x 12
		8'd22, 	 // 2 x 11
		8'd20, 	 // 2 x 10
		8'd18, 	 // 2 x 9
		8'd16, 	 // 2 x 8
		8'd14, 	 // 2 x 7
		8'd12, 	 // 2 x 6
		8'd10, 	 // 2 x 5
		8'd8, 	 // 2 x 4
		8'd6, 	 // 2 x 3
		8'd4, 	 // 2 x 2
		8'd2, 	 // 2 x 1
		8'd0, 	 // 2 x 0
		8'd15, 	 // 1 x 15
		8'd14, 	 // 1 x 14
		8'd13, 	 // 1 x 13
		8'd12, 	 // 1 x 12
		8'd11, 	 // 1 x 11
		8'd10, 	 // 1 x 10
		8'd9, 	 // 1 x 9
		8'd8, 	 // 1 x 8
		8'd7, 	 // 1 x 7
		8'd6, 	 // 1 x 6
		8'd5, 	 // 1 x 5
		8'd4, 	 // 1 x 4
		8'd3, 	 // 1 x 3
		8'd2, 	 // 1 x 2
		8'd1, 	 // 1 x 1
		8'd0, 	 // 1 x 0
		8'd0, 	 // 0 x 15
		8'd0, 	 // 0 x 14
		8'd0, 	 // 0 x 13
		8'd0, 	 // 0 x 12
		8'd0, 	 // 0 x 11
		8'd0, 	 // 0 x 10
		8'd0, 	 // 0 x 9
		8'd0, 	 // 0 x 8
		8'd0, 	 // 0 x 7
		8'd0, 	 // 0 x 6
		8'd0, 	 // 0 x 5
		8'd0, 	 // 0 x 4
		8'd0, 	 // 0 x 3
		8'd0, 	 // 0 x 2
		8'd0, 	 // 0 x 1
		8'd0	 	 // 0 x 0
};

mult =  ROM[{address1, address2}];
endfunction
